library IEEE;
use IEEE.STD_LOGIC_1164.all;

package TOP_PACKAGE is

-- type <new_type> is
--  record
--    <type_name>        : std_logic_vector( 7 downto 0);
--    <type_name>        : std_logic;
-- end record;
--
-- Declare constants
--
-- constant <constant_name>		: time := <time_unit> ns;
-- constant <constant_name>		: integer := <value;
--
-- Declare functions and procedure
--
-- function <function_name>  (signal <signal_name> : in <type_declaration>) return <type_declaration>;
-- procedure <procedure_name> (<type_declaration> <constant_name>	: in <type_declaration>);
--
	CONSTANT LW : STD_LOGIC_VECTOR(6 DOWNTO 0):= "0000011";
	CONSTANT SW : STD_LOGIC_VECTOR(6 DOWNTO 0):= "0100011";
	CONSTANT BEQ : STD_LOGIC_VECTOR(6 DOWNTO 0):= "1100111";
	CONSTANT R : STD_LOGIC_VECTOR(6 DOWNTO 0):= "0110011";
	

end TOP_PACKAGE;

package body TOP_PACKAGE is

---- Example 1
--  function <function_name>  (signal <signal_name> : in <type_declaration>  ) return <type_declaration> is
--    variable <variable_name>     : <type_declaration>;
--  begin
--    <variable_name> := <signal_name> xor <signal_name>;
--    return <variable_name>; 
--  end <function_name>;

---- Example 2
--  function <function_name>  (signal <signal_name> : in <type_declaration>;
--                         signal <signal_name>   : in <type_declaration>  ) return <type_declaration> is
--  begin
--    if (<signal_name> = '1') then
--      return <signal_name>;
--    else
--      return 'Z';
--    end if;
--  end <function_name>;

---- Procedure Example
--  procedure <procedure_name>  (<type_declaration> <constant_name>  : in <type_declaration>) is
--    
--  begin
--    
--  end <procedure_name>;


 
end TOP_PACKAGE;
